// mips_decode: a decoder for MIPS arithmetic instructions
//
// alu_op       (output) - control signal to be sent to the ALU
// writeenable  (output) - should a new value be captured by the register file
// rd_src       (output) - should the destination register be rd (0) or rt (1)
// alu_src2     (output) - should the 2nd ALU source be a register (0) or an immediate (1)
// except       (output) - set to 1 when we don't recognize an opdcode & funct combination
// control_type (output) - 00 = fallthrough, 01 = branch_target, 10 = jump_target, 11 = jump_register 
// mem_read     (output) - the register value written is coming from the memory
// word_we      (output) - we're writing a word's worth of data
// byte_we      (output) - we're only writing a byte's worth of data
// byte_load    (output) - we're doing a byte load
// lui          (output) - the instruction is a lui
// slt          (output) - the instruction is an slt
// addm         (output) - the instruction is an addm
// opcode        (input) - the opcode field from the instruction
// funct         (input) - the function field from the instruction
// zero          (input) - from the ALU
//

module mips_decode(alu_op, writeenable, rd_src, alu_src2, except, control_type,
                   mem_read, word_we, byte_we, byte_load, lui, slt, addm,
                   opcode, funct, zero);
    output [2:0] alu_op;
    output       writeenable, rd_src, alu_src2, except;
    output [1:0] control_type;
    output       mem_read, word_we, byte_we, byte_load, lui, slt, addm;
    input  [5:0] opcode, funct;
    input        zero;
	wire beq, bne, j, jr, lw, lbu, sw, sb;
	wire w1, addi, andi, ori, xori, add, sub, and1, or1, nor1, xor1;


	assign w1 = (opcode == 6'b0);
	assign addi = (opcode == 6'b1000);
	assign andi = (opcode == 6'b1100);
	assign ori = (opcode == 6'b1101);
	assign xori = (opcode == 6'b1110);
	assign add = w1 & (funct == 6'b100000);
	assign sub = w1 & (funct == 6'b100010);
	assign and1 = w1 & (funct == 6'b100100);
	assign or1 = w1 & (funct == 6'b100101);
	assign nor1 = w1 & (funct == 6'b100111);
	assign xor1 = w1 & (funct == 6'b100110);

	assign beq = (opcode == `OP_BEQ);
	assign j = (opcode == `OP_J);
	assign bne = (opcode == `OP_BNE);
	assign jr = w1 &  (funct == `OP0_JR);
	assign lw = (opcode == `OP_LW);
	assign lbu = (opcode == `OP_LBU);
	assign sw = (opcode == `OP_SW);
	assign sb = (opcode == `OP_SB);
	assign addm = w1 & (funct == `OP0_ADDM);



	assign lui = (opcode == 6'b001111);
	assign slt = w1 & (funct == 6'b101010);
	assign rd_src = addi|andi|ori|xori|lbu|lui|lw;
	assign alu_src2 = addi|andi|ori|xori|lw|lbu|sw|sb;
	assign mem_read = (lw|lbu|addm); 
	assign word_we = sw; 
	assign byte_we = sb;
	assign byte_load = lbu;
	

	assign control_type[0] = ((beq& zero)|(bne& ~zero)|jr);
	assign control_type[1] = j|jr;
	assign alu_op[0] = sub|or1|xor1|ori|xori|beq|bne|slt;
	assign alu_op[1] = addi|xori|add|sub|nor1|xor1|beq|bne|sb|sw|lw|lbu|slt|addm;
	assign alu_op[2] = andi|ori|xori|and1|or1|nor1|xor1;
	assign writeenable = add|sub|and1|or1|nor1|xor1|addi|andi|ori|xori|lbu|lui|lw|slt|addm;
	assign except = ~(add|sub|and1|or1|nor1|xor1|addi|andi|ori|xori|lbu|lui|lw|slt|j|jr|sw|sb|bne|beq|addm);	

	
endmodule // mips_decode

